// SPDX-FileCopyrightText: © 2020-2024 The Bluespec Authors
// SPDX-License-Identifier: BSD-3-Clause

`include "bluespec.svh"

// -- AMALGAMATE: start --
// ---------------------------------------------------------------------------------------------------------------------

// __BSC_NULL__: An empty module to be used as a placeholder.
module __BSC_NULL__ (); endmodule: __BSC_NULL__ // # MARK: __BSC_NULL__

// ---------------------------------------------------------------------------------------------------------------------

`ifdef __BSC_SHIM_V1_PRIMS__
module BypassWire0 (); endmodule
`endif // __BSC_SHIM_V1_PRIMS__

// ---------------------------------------------------------------------------------------------------------------------
// -- AMALGAMATE: end --
